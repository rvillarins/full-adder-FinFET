*Full adder 

* Libraries
.include 16nm_PTM_HP.pm

* Transistor's W parameters (tenologies)

.param wp=32n
.param wn=16n
.param supply = 0.7

* VDD and power suplies
VVdd    VDD gnd supply
.global VDD

Va   A   gnd pwl(0 0 1n 0           2n 0           3n 0 3.01n 0.7 4n 0.7         5n 0.7         6n 0.7 6.01n 0 7n 0 7.01n 0.7 8n 0.7 8.01n 0 9n 0           10n 0            11n 0              12n 0            13n 0            14n 0            15n 0              16n 0   16.01n 0.7 17n 0.7 17.01n 0 18n 0   18.01n 0.7 19n 0.7          20n 0.7          21n 0.7 21.01n 0   22n 0            23n 0            24n 0)
Vb   B   gnd pwl(0 0 1n 0           2n 0 		   3n 0 3.01n 0.7 4n 0.7         5n 0.7         6n 0.7 6.01n 0 7n 0           8n 0           9n 0 9.01n 0.7 10n 0.7 10.01n 0 11n 0   11.01n 0.7 12n 0.7 12.01n 0 13n 0 13.01n 0.7 14n 0.7 14.01n 0 15n 0   15.01n 0.7 16n 0.7            17n 0.7          18n 0.7 18.01n 0   19n 0            20n 0            21n 0   21.01n 0.7 22n 0.7          23n 0.7          24n 0.7)
VCin CIN gnd pwl(0 0 1n 0 1.01n 0.7 2n 0.7 2.01n 0 3n 0           4n 0 4.01n 0.7 5n 0.7 5.01n 0 6n 0           7n 0           8n 0           9n 0 9.01n 0.7 10n 0.7          11n 0.7            12n 0.7          13n 0.7          14n 0.7          15n 0.7 15.01n 0   16n 0              17n 0            18n 0              19n 0 19.01n 0.7 20n 0.7 20.01n 0 21n 0              22n 0 22.01n 0.7 23n 0.7 23.01n 0 24n 0)     
                                                                                                                                                                             
**************************************Circuito************************************* 
***********************************Subcircuito Nand********************************
.subckt NAND A B OUT
MP1 VDD a out VDD PMOS w=wp l=16n 
MP2 VDD b out VDD PMOS w=wp l=16n

MN1 out a N1  gnd NMOS w=wn l=16n 
MN2 N1  b gnd gnd NMOS w=wn l=16n
.ends NAND

***********Somador projetado a partir de portas lógicas NAND de 2 entradas*********
X1 A   B  N2   NAND
X2 A   N2 N4   NAND
X3 N2  B  N3   NAND
X4 N4  N3 N5   NAND
X5 CIN N5 N6   NAND
X6 CIN N6 N7   NAND
X7 N5  N6 N8   NAND
X8 N6  N2 COUT NAND
X9 N7  N8 SUM  NAND

*************************************Capacitores************************************
Ccout COUT gnd 1f
Csum  SUM  gnd 1f

**********************************Tipo de simulação*********************************
.TRAN 0.01n 24n

*****Medições de Atraso em relação as saidas de Soma e Carry-out do somador*********
.MEASURE TRAN td_lh_c0 TRIG     v(CIN) VAL=0.35 RISE=1 TARG v(SUM) VAL=0.35 RISE=1
.MEASURE TRAN td_hl_c0 TRIG     v(CIN) VAL=0.35 FALL=1 TARG v(SUM) VAL=0.35 FALL=1
							    
.MEASURE TRAN td_lh_c1 TRIG     v(CIN) VAL=0.35 RISE=2 TARG v(SUM) VAL=0.35 RISE=2
.MEASURE TRAN td_hl_c1 TRIG     v(CIN) VAL=0.35 FALL=2 TARG v(SUM) VAL=0.35 FALL=2
							    
.MEASURE TRAN td_lh_a0 TRIG     v(A)   VAL=0.35 RISE=2 TARG v(SUM) VAL=0.35 FALL=3
.MEASURE TRAN td_hl_a0 TRIG     v(A)   VAL=0.35 FALL=2 TARG v(SUM) VAL=0.35 FALL=3
							    
.MEASURE TRAN td_lh_b0 TRIG     v(B)   VAL=0.35 FALL=2 TARG v(SUM) VAL=0.35 RISE=4
.MEASURE TRAN td_hl_c0 TRIG     v(B)   VAL=0.35 RISE=3 TARG v(SUM) VAL=0.35 FALL=4

.MEASURE TRAN td_lh_bcout0 TRIG v(B)   VAL=0.35 RISE=3 TARG v(COUT) VAL=0.35 RISE=5
.MEASURE TRAN td_hl_bcout0 TRIG v(B)   VAL=0.35 FALL=3 TARG v(COUT) VAL=0.35 FALL=5
									   
.MEASURE TRAN td_lh_acout0 TRIG v(A)   VAL=0.35 RISE=3 TARG v(COUT) VAL=0.35 RISE=6
.MEASURE TRAN td_hl_acout0 TRIG v(A)   VAL=0.35 FALL=3 TARG v(COUT) VAL=0.35 FALL=6

.MEASURE TRAN td_lh_ccout0 TRIG v(CIN) VAL=0.35 RISE=4 TARG v(COUT) VAL=0.35 RISE=7
.MEASURE TRAN td_hl_ccout0 TRIG v(CIN) VAL=0.35 FALL=4 TARG v(COUT) VAL=0.35 FALL=7

.MEASURE TRAN td_lh_ccout1 TRIG v(CIN) VAL=0.35 RISE=5 TARG v(COUT) VAL=0.35 RISE=8
.MEASURE TRAN td_hl_ccout1 TRIG v(CIN) VAL=0.35 FALL=5 TARG v(COUT) VAL=0.35 FALL=8

****************************Medição de energia e Potencia***************************
.measure tran energ_FAvdd INTEG i(vvdd) from=0.01n to=24n
.measure tran energ_FAva  INTEG i(vva)  from=0.01n to=24n
.measure tran energ_FAvb  INTEG i(vvb)  from=0.01n to=24n
.measure tran energ_FAvc  INTEG i(vvc)  from=0.01n to=24n


.measure tran avgi_a   AVG i(va)   from=0.01n to=24n 
.measure tran avgi_b   AVG i(vb)   from=0.01n to=24n 
.measure tran avgi_cin AVG i(vcin) from=0.01n to=24n 

.measure tran powera PARAM = ((((avgi_a)) + (avgi_b * (-1)) + (avgi_cin)) * 0.7)

.control
set color0=magenta
set xbrushwidth=3
run
display 
*plot v(A)
*plot v(B)
*plot v(CIN)
*plot v(COUT)
*plot v(SUM)
.endc

.end